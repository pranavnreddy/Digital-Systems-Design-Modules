// Code your testbench here
// or browse Examples
`include "lab2_3_tb.sv"