// Code your testbench here
// or browse Examples
//`include "lab2_2_tb.sv"
`include "lab2_tb_file.sv"
