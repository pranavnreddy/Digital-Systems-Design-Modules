// Code your design here
`include "robsmult.sv"
`include "addsub.sv"
`include "robs_control_unit_micro.sv"
`include "robs_data_path.sv"
`include "counter_down.sv"
`include "mux2.sv"
`include "mux5.sv"
`include "mux3.sv"
`include "register_hl.sv"
`include "register.sv"
`include "rom.sv"
`include "upc_reg.sv"
`include "right_shift_register.sv"