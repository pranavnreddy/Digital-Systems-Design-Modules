// Code your testbench here
// or browse Examples
`include "robertsonstest.sv"