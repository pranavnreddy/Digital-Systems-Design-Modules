// Code your design here
`include "alarm.sv"
`include "ct_mod_N.sv"
`include "lcd_int3.sv"
`include "struct_diag.sv"